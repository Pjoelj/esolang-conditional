rstv r0 0
rstr r1 r0
radr r0 r1