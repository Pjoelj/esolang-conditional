vwtm 72 0
vwtm 101 1
vwtm 108 2
vwtm 108 3
vwtm 111 4
vwtm 44 5
vwtm 32 6
vwtm 87 7
vwtm 111 8
vwtm 114 9
vwtm 108 10
vwtm 100 11
vwtm 33 12
vwtm 10 13
moup 0 14